** Profile: "SCHEMATIC1-a"  [ C:\Users\DTIC\Desktop\P1_Pspice\P1_Pspice-PSpiceFiles\SCHEMATIC1\a.sim ] 

** Creating circuit file "a.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../librarii/smls14bet.lib" 
* From [PSPICE NETLIST] section of C:\Users\DTIC\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 2ms 0 50ns 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
