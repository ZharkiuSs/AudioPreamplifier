** Profile: "SCHEMATIC1-AmplificareMin"  [ C:\Users\Eduard\Desktop\P1Eu\P1_2024_432B_Gherghel_Eduard-Mihai_PaCT_N5_CISLite\SCHEMATIC\P1_PspiceVechi\P1_Pspice-PSpiceFiles\SCHEMATIC1\AmplificareMin.sim ] 

** Creating circuit file "AmplificareMin.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../librarii/smls14bet.lib" 
* From [PSPICE NETLIST] section of C:\Users\Eduard\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 4ms 0 50ns 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
